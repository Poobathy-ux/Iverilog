module and_gate_p (c,a,b);
output wire c;
 input wire a,b;
and aq(c,a,b);
endmodule   
            
